library verilog;
use verilog.vl_types.all;
entity testbench_alu is
end testbench_alu;
