module testbench_prog();
// Declare inputs as regs and outputs as wires
reg clk;
 wire	taken;
 wire	halt;
 wire	[3:0] alu_NZCV;
 wire	[7:0] alu_reg1;
 wire	[7:0] alu_reg2;
 wire	[7:0] alu_result;
 wire	[8:0] instr_out;
 wire	[7:0] mem_addr;
 wire	[7:0] mem_datain;
 wire	[7:0] mem_out;
 wire	[7:0] pc;
 wire	[7:0] reg_in;
 wire	[1:0] reg_in_src;
 wire	[7:0] reg_out1;
 wire	[7:0] reg_out2;
 wire	[2:0] special_func;
wire	[3:0] dec_full;
wire	[7:0] dec_imm;
wire	[7:0] dec_imm_br;
wire	[2:0] dec_r1;
wire	[2:0] dec_r2;
wire	con_spec_op;
wire	con_write_reg;
wire	con_read_reg;
wire	reg_ldst;
wire	[1:0] reg_aro;
wire	[2:0] dec_rw;
wire	branch;
wire	[7:0] target_pc;
wire	[7:0] new_pc;
wire	[15:0] dyn;
wire	[2:0] pipe_state;

// Initialize all variables
// Clock generator
initial begin
clk=0;
end
always begin
#5 clk = ~clk; // Toggle clock every 5 ticks
// this makes the clock cycle 10 ticks
end
// the following creates an instance of our program_counter register.

// I copied this code verbatim from the pc_schematic.v that was
// generated by Quartus when I created the .v file from the .bdf.

 pc_schematic pc_schem_inst(
	.clk(clk),
	.taken(taken),
	.halt(halt),
	.alu_NZCV(alu_NZCV),
	.alu_reg1(alu_reg1),
	.alu_reg2(alu_reg2),
	.alu_result(alu_result),
	.instr_out(instr_out),
	.pc(pc),
	.mem_addr(mem_addr),
	.mem_datain(mem_datain),
	.mem_out(mem_out),
	.reg_in(reg_in),
	.reg_in_src(reg_in_src),
	.reg_out1(reg_out1),
	.reg_out2(reg_out2),
	.special_func(special_func),
	.dec_full(dec_full),
	.dec_imm(dec_imm),
	.dec_imm_br(dec_imm_br),
	.dec_r1(dec_r1),
	.dec_r2(dec_r2),
	.con_spec_op(con_spec_op),
	.con_write_reg(con_write_reg),
	.con_read_reg(con_read_reg),
	.reg_ldst(reg_ldst),
	.reg_aro(reg_aro),
	.dec_rw(dec_rw),
	.branch(branch),
	.target_pc(target_pc),
	.new_pc(new_pc),
	.dyn(dyn),
	.pipe_state(pipe_state)
);
	
endmodule