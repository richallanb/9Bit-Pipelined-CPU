library verilog;
use verilog.vl_types.all;
entity testbench_prog is
end testbench_prog;
