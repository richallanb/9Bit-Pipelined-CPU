module testbench_alu();
// Declare inputs as regs and outputs as wires
reg clk;
reg [1:0] aro;
reg spec;
reg [2:0]spec_fun;
reg [7:0]r1;
reg [7:0]r2;
reg [7:0]r3;
reg [7:0]r4;
reg ALon;

wire [7:0] res;
wire [3:0] NZCV;
// Initialize all variables
initial begin
clk = 1; // initial value of clock
ALon = 0; // initial value of ALUon
spec = 0; // initial value of special_op (off)
spec_fun = 3'b000; // initial value of special function
aro = 2'b00; // initial value of aro (add)
#10 r1 = 8'd3;
#10 r2 = 8'd5;
#10 // wait a cycle, make sure result wasn't computed
#10 ALon = 1; r1=8'd5; r2=8'd1; // set ALon high  -> 5+1
#10 aro=2'b01; r1=8'd5; r2=8'd1;// 5-1
#10 r1=8'd5; r2=8'd5;// 5-5
#10 r1=8'd3; r2=8'd6;// 3-6
#10 aro=2'b10; r1=8'd5; r2=8'd5; // cmp 5,5
#10 r1=8'd6; r2=8'd2; // cmp 6,2
#10 r1=8'd4; r2=8'd10; // cmp 4,10
#10 aro=2'b11; r1=8'd5; r2=8'd5; // slt 5,5
#10 r1=8'd6; r2=8'd2; // slt 6,2
#10 r1=8'd4; r2=8'd10; // slt 4,10
#10 r1=8'd0; r2=8'd255; // slt 4,10
#10 spec=1; spec_fun =3'b000; r1=0; r2=3; r3=2; r4=0; // MFL
#10 spec_fun =3'b001; r1=0; r2=8'b10111110; // SPC
#10 spec_fun =3'b001; r1=1; r2=8'b11110010; // SPC
#10 spec_fun =3'b001; r1=2; r2=8'b10110110; // SPC
#10 spec_fun =3'b010; r1=0; r2=3; r3=2; r4=0; // MFH
#10 spec_fun =3'b011; r1=3; r2=8; // ISC
#10 spec_fun =3'b100; r1=10; // INC
#10 spec_fun =3'b101; r1=107; // SM



end
// Clock generator
always begin
#5 clk = ~clk; // Toggle clock every 5 ticks
// this makes the clock cycle 10 ticks
end
// the following creates an instance of our program_counter register.

// I copied this code verbatim from the pc_schematic.v that was
// generated by Quartus when I created the .v file from the .bdf.
alu alu_inst(
.aro(aro),
.special_op(spec),
.special_func(spec_fun),
.reg1(r1),
.reg2(r2),
.reg3(r3),
.reg4(r4),
.ALUon(ALon),
.clk(clk),
.result(res),
.NZCV(NZCV));
endmodule