library verilog;
use verilog.vl_types.all;
entity testbench_reg is
end testbench_reg;
