module testbench();
// Declare inputs as regs and outputs as wires
reg clk;
reg wenable;
reg reset;
reg start;
reg branch;
reg taken;
reg [7:0]target;
wire [7:0] currentpc;
wire [7:0] newpc;
wire [8:0] instr;
// Initialize all variables
initial begin
clk = 1; // initial value of clock
reset = 0; // initial value of reset
wenable = 0; // initial value of wenable
#10 reset = 1; // use reset to set pc to 0
#10 reset = 0; // end of reset pulse.
#10 // wait a cycle, make sure the PC doesn't change
#10 wenable = 1; start=1;
#10 // wait a cycle, pc should increment to 1
#10 // cycle pc = 2
#10 branch = 1; taken=1; target=7;//pc should go to 7
#10 branch = 0;
#10 //pc should be 9
#10 //pc should be 10
#10 start = 0;
#10 //pc should keep its value
#10 //pc should keep its value
#10 branch = 1; taken=0;
#10 //nothing should change
#10 target = 8'b0000110;
#10 start = 1; //pc should now be set to 11 (branch not taken)
#10 start = 0; //stop pc
#10 reset = 1; //see if reset works when wenable high
#10 reset = 0; wenable = 0;
end
// Clock generator
always begin
#5 clk = ~clk; // Toggle clock every 5 ticks
// this makes the clock cycle 10 ticks
end
// the following creates an instance of our program_counter register.

// I copied this code verbatim from the pc_schematic.v that was
// generated by Quartus when I created the .v file from the .bdf.
program_counter b2v_inst(
.clock(clk),
.wenable_i(wenable),
.reset_i(reset),
.newpc_i(newpc),
.pc_o(currentpc));

next_pc_logic fetch_inst(
.start(start),
.currentpc(currentpc),
.branch(branch),
.target(target),
.taken(taken),
.clk(clk),
.pc_o(newpc));

instruction_rom instr_rom(.clk(clk), .pc_line(newpc), .instr_out(instr));

endmodule